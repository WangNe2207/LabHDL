library verilog;
use verilog.vl_types.all;
entity tb_add is
end tb_add;
